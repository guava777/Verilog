module hello;
    initial begin
        $display("Hello");
        $finish;
    end

endmodule